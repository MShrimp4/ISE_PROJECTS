`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:53:33 05/03/2019 
// Design Name: 
// Module Name:    gt_board 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module gt_board(
	input wire [3:0] a;
	input wire [3:0] b;
	output wire agtb;
    );
	

endmodule
